library verilog;
use verilog.vl_types.all;
entity TestbenchControlUnit is
end TestbenchControlUnit;
